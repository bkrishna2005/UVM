class dff_driver extends uvm_driver#(dff_transaction)
  `uvm_component_utils(dff_driver)
  
endclass